
`define OPCODE_ALU  7'b0110011
`define OPCODE_LOAD 7'b0000011
`define OPCODE_LOAD_IMM 7'b0000011